netcdf ssat {
dimensions:
  dim = 2 ;
  n = 11 ;
  nlayer = 4 ;
  nparam = 10 ;
variables:
  double elevation_profile(dim, n) ;
    elevation_profile:units = "feet" ;
  double stratum(nlayer, nparam) ;
data:
 elevation_profile = 0.0, 15.0, 15.0, 15.0, 39.0, -2.6, 45.0, -2.6, 84.5,
   -31.8, 108.0, -31.8, 133.3, -31.8, 165.0, -2.6, 195.0, -2.6, 218.0, 15.0,
   225.0, 15.0, 0.00
     4
   4.0  17.28  30.00   0.00   0.00   0.00   0.00   0.00   0.00   0.00
 -10.0  20.75   0.00  50.77   0.21   0.00   0.00   0.00   0.00   0.00
 -30.0  20.11   0.00  29.69   0.24   0.00   0.00   0.00   0.00   0.00
 -40.0  20.11   0.00  37.36   0.26   0.00   0.00   0.00   0.00   0.00
     0
