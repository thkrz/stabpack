netcdf pwp {
dimensions:
  m = 2 ;
  n = 2 ;
variables:
  float map(m, n) ;
    map:dx = 1.0 ;
    map:dy = 1.0 ;
    map:origin_x = 0.0 ;
    map:origin_y = 0.0 ;
  :title = "Pore water pressure" ;
data:
  map =
  1, 2, NaN, 4 ;
}
